module t_file();
    



endmodule